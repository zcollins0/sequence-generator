* SPICE3 file created from NOR2X1.ext - technology: scmos
.include ~/model_t36s.sp
.option scale=0.3u
.param vdd=5V

vdd vdd 0 vdd

Va a 0 PWL(0 0 10n 0 20n 0 20.1n 5V 40n 5V 40.1n 0V)
Vb b 0 PWL(0 0 10n 0 10.1n 5V 30n 5V 30.1n 0V)
.options post=2
.tran 1p 50n

M1000 a_9_54# a vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=200 ps=90
M1001 y b a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1002 y a gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=100 ps=60
M1003 gnd b y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
C0 gnd Gnd 2.71fF
C1 vdd Gnd 8.40fF
