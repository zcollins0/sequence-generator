magic
tech scmos
timestamp 1072202993
<< polysilicon >>
rect 0 0 150 2900
<< end >>
