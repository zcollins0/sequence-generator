* SPICE3 file created from AND2X1.ext - technology: scmos

.include ~/model_t36s.sp
.option scale=0.3u
.param vdd=5V

VA A 0 PWL(0 0V 10n 0V 10.1n 5V 20n 5V 20.1n 0V 50n 0V)
VB B 0 PWL(0 0V 10n 0V 10.1n 5V 20n 5V 50n 5V)

.options post=2
.tran 1p 50n

vdd vdd 0 vdd
M1000 a_2_6# A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=220 ps=102
M1001 vdd B a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 Y a_2_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1003 a_9_6# A a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M1004 gnd B a_9_6# Gnd nfet w=20 l=2
+  ad=110 pd=52 as=0 ps=0
M1005 Y a_2_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
C0 Y Gnd 2.26fF
C1 gnd Gnd 2.81fF
C2 a_2_6# Gnd 2.24fF
C3 vdd Gnd 10.25fF
