* SPICE3 file created from NOR2X1.ext - technology: scmos

.option scale=0.3u

M1000 a_9_54# a vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=200 ps=90
M1001 y b a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1002 y a gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=100 ps=60
M1003 gnd b y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
C0 gnd Gnd 2.71fF
C1 vdd Gnd 8.40fF
