* SPICE3 file created from TBUFX1.ext - technology: scmos
.include ~/model_t36s.sp
.option scale=0.3u
.param vdd=5V

vdd vdd 0 vdd
VEN en 0 PWL(0 5V)
VD a 0 PWL(0 0 10n 0 10.1n 5V 25n 5V 25.1n 0V)
.options post=2
.tran 1p 50n

M1000 a_9_6# en vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=300 ps=140
M1001 a_26_54# a_9_6# Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=200 ps=90
M1002 vdd a a_26_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 a_9_6# en gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=150 ps=80
M1004 a_26_6# en Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M1005 gnd a a_26_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
C0 a_9_6# vdd 2.08fF
C1 gnd Gnd 3.85fF
C2 a_9_6# Gnd 2.38fF
C3 vdd Gnd 9.98fF
