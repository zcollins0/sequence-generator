magic
tech scmos
timestamp 1541537479
<< nwell >>
rect -8 48 40 105
<< ntransistor >>
rect 7 6 9 26
rect 12 6 14 26
rect 20 6 22 16
<< ptransistor >>
rect 7 74 9 94
rect 15 74 17 94
rect 23 74 25 94
<< ndiffusion >>
rect 6 6 7 26
rect 9 6 12 26
rect 14 6 15 26
rect 19 6 20 16
rect 22 6 23 16
<< pdiffusion >>
rect 6 74 7 94
rect 9 74 10 94
rect 14 74 15 94
rect 17 74 18 94
rect 22 74 23 94
rect 25 74 26 94
<< ndcontact >>
rect 2 6 6 26
rect 15 6 19 26
rect 23 6 27 16
<< pdcontact >>
rect 2 74 6 94
rect 10 74 14 94
rect 18 74 22 94
rect 26 74 30 94
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 23 94 25 96
rect 7 41 9 74
rect 15 53 17 74
rect 6 37 9 41
rect 15 39 17 49
rect 7 26 9 37
rect 12 37 17 39
rect 12 26 14 37
rect 23 33 25 74
rect 24 30 25 33
rect 20 16 22 29
rect 7 4 9 6
rect 12 4 14 6
rect 20 4 22 6
<< polycontact >>
rect 13 49 17 53
rect 2 37 6 41
rect 20 29 24 33
<< metal1 >>
rect 7 103 11 111
rect -2 102 34 103
rect 2 98 14 102
rect 18 98 34 102
rect -2 97 34 98
rect 2 94 6 97
rect 18 94 22 97
rect 11 71 14 74
rect 11 68 23 71
rect 6 53 17 57
rect -2 33 6 37
rect 20 33 23 68
rect 27 43 30 74
rect 27 39 34 43
rect 9 30 20 33
rect 9 29 12 30
rect 3 26 12 29
rect 27 19 30 39
rect 23 16 30 19
rect 15 3 19 6
rect -2 2 34 3
rect 2 -2 14 2
rect 18 -2 34 2
rect -2 -3 34 -2
rect 6 -7 10 -3
<< m1p >>
rect 26 63 30 67
rect 10 53 14 57
rect 2 33 6 37
<< labels >>
rlabel m1p 28 65 28 65 6 Y
rlabel m1p 12 55 12 55 6 B
rlabel metal1 4 100 4 100 6 vdd
rlabel metal1 4 0 4 0 8 gnd
rlabel m1p 4 35 4 35 6 A
rlabel metal1 7 107 11 111 5 Vdd
rlabel metal1 30 39 34 43 1 Y
rlabel metal1 -2 33 2 37 1 A
rlabel metal1 6 -7 10 -3 1 Gnd
rlabel metal1 6 53 10 57 1 B
<< end >>
